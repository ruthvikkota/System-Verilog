class transaction;
  rand bit a, b;
  bit sum, carry;
endclass

