interface intf;
logic a,b;
logic d0,d1,d2,d3;
endinterface

