class transaction;
rand bit a,b;
bit d0,d1,d2,d3;
endclass

